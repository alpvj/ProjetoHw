module Controle(input logic overflow, DIV0, clk, EQF, GTF, input logic [5:0] OpCode, funct,
output logic PCWrite, MemCtrl, IRWrite, A_Control, B_Control, RegControl, ALUOutControl, EPCWrite, MDControl, HI_Control, LO_Control,
output logic [1:0] IorD, ALUSrcA, ALUSrcB, ExcpCtrl, ShiftSrc, ShiftAmt, SSControl, LSControl,
output logic [2:0] RegDst, PCSource, ALUControl, ShiftControl,
output logic [3:0] DataSrc,
output logic [6:0] estado,
output logic reset);//11 + 8 + 4 + 1 = 24 sinais de controle

/*
PCWrite = 1'b0;
MemCtrl = 1'b0;
IRWrite = 1'b0;
A_Control = 1'b0;
B_Control = 1'b0;
RegControl = 1'b0;
ALUOutControl = 1'b0;
EPCWrite = 1'b0;
MDControl = 1'b0;
HI_Control = 1'b0;
LO_Control = 1'b0;
IorD = 2'b00;
ALUSrcA = 2'b00;
ALUSrcB = 2'b00;
ExcpCtrl = 2'b00;
ShiftSrc = 2'b00;
ShiftAmt = 2'b00;
SSControl = 2'b00;
LSControl = 2'b00;
RegDst = 3'b000;
PCSource = 3'b000;
ALUControl = 3'b000;
ShiftControl = 3'b000;
DataSrc = 4'b0000;
estado = 7'b0000000;
*/

//Estados
parameter Fetch1 = 7'd0;
parameter Espera1Fetch = 7'd1;
parameter Espera2Fetch = 7'd2;
parameter Fetch2 = 7'd3;
parameter Decode1 = 7'd4;
parameter EsperaDecode = 7'd5;
parameter Decode2 = 7'd6;
parameter Instrucao = 7'd7;

parameter Add2 = 7'd8;
parameter Sub2 = 7'd9;
parameter And2 = 7'd10;
parameter AddSubAnd = 7'd11;
parameter AddSubAnd2 = 7'd12;
parameter Addi2 = 7'd13;
parameter Addi3 = 7'd14;
parameter Addi4 = 7'd15;
parameter Break2 = 7'd16;
parameter Break3 = 7'd17;
parameter Rte2 = 7'd18;
parameter Sll2 = 7'd19;
parameter Sll3 = 7'd20;
parameter Sll4 = 7'd21;
parameter Sllv2 = 7'd22;
parameter Sllv3 = 7'd23;
parameter Srl2 = 7'd24;
parameter Srl3 = 7'd25;
parameter Sra2 = 7'd26;
parameter Sra3 = 7'd27;
parameter Srav2 = 7'd28;
parameter Srav3 = 7'd29;
parameter Addiu2 = 7'd30;
parameter Addiu3 = 7'd31;
parameter Slt2 = 7'd32;
parameter Slt3 = 7'd33;
parameter jr2 = 7'd34;
parameter xchg2 = 7'd35;
parameter xchg3 = 7'd36;
parameter xchg4 = 7'd37;
parameter j2 = 7'd38;
parameter jal2 = 7'd39;
parameter lui2 = 7'd40;
parameter lui3 = 7'd41;
parameter lui4 = 7'd42;
parameter slti2 = 7'd43;
parameter slti3 = 7'd44;
parameter beq2 = 7'd45;
parameter beq3 = 7'd46;
parameter beq4 = 7'd47;
parameter bne2 = 7'd48;
parameter bne3 = 7'd49;
parameter ble2 = 7'd50;
parameter ble3 = 7'd51;
parameter bgt2 = 7'd52;
parameter bgt3 = 7'd53;
parameter OVERFLOW = 7'd54;
parameter sb2 = 7'd55;
parameter sb3 = 7'd56;
parameter sbWait = 7'd57;
parameter sbWait2 = 7'd58;
parameter lb2 = 7'd59;
parameter lb3 = 7'd60;
parameter lbWait = 7'd61;
parameter lbWait2 = 7'd62;
parameter lbWait3 = 7'd63;
parameter lh2 = 7'd64;
parameter lh3 = 7'd65;
parameter lhWait = 7'd66;
parameter lhWait2 = 7'd67;
parameter lhWait3 = 7'd68;
parameter lw2 = 7'd69;
parameter lw3 = 7'd70;
parameter lwWait = 7'd71;
parameter lwWait2 = 7'd72;
parameter lwWait3 = 7'd73;
parameter sh2 = 7'd74;
parameter sh3 = 7'd75;
parameter shWait = 7'd76;
parameter shWait2 = 7'd77;
parameter sw2 = 7'd78;
parameter sw3 = 7'd79;
parameter swWait = 7'd80;
parameter swWait2 = 7'd81;
parameter blm2 = 7'd82;
parameter blm3 = 7'd83;
parameter blm4 = 7'd84;
parameter blm5 = 7'd85;
parameter blm6 = 7'd86;
parameter overflow2 = 7'd86;
parameter overflow3 = 7'd87;
parameter overflow4 = 7'd88;
parameter overflow5 = 7'd89;
parameter INEXISTENTE = 7'd90;
parameter inexistente2 = 7'd91;
parameter inexistente3 = 7'd92;
parameter inexistente4 = 7'd93;
parameter inexistente5 = 7'd94;


//Func do Tipo R
parameter ADD = 6'b100000;//done
parameter SUB = 6'b100010;//done
parameter AND = 6'b100100;//done
parameter BREAK = 6'b001101;//done
parameter RTE = 6'b010011;//done
parameter SLL = 6'b000000;//done
parameter SLLV = 6'b000100;//done
parameter SRA = 6'b000011;//done
parameter SRAV = 6'b000111;//done
parameter SRL = 6'b000010;//done
parameter SLT = 6'b101010;//done
parameter JR = 6'b001000;//done
parameter XCHG = 6'b000101;//done


//Opcodes
parameter ARIT = 6'b000000;
//Tipo I
parameter ADDI = 6'b001000;
parameter ADDIU = 6'b001001;//done
parameter LUI = 6'b001111;//done
parameter SLTI = 6'b001010;//done
parameter BEQ = 6'b000100;//done
parameter BNE = 6'b000101;//done
parameter BLE = 6'b000110;//done
parameter BGT = 6'b000111;//done
parameter LB = 6'b100000;//done
parameter LH = 6'b100001;//done
parameter LW = 6'b100011;//done
parameter SB = 6'b101000;//done
parameter SH = 6'b101001;//done
parameter SW = 6'b101011;//done
parameter BLM = 6'b000001;//done
//Func do Tipo J
parameter J = 6'b000010;//done
parameter JAL = 6'b000011;//done



initial begin
	estado = Fetch1;
	reset = 1'b1;
end

always @(posedge clk) begin
	if (reset) begin
		reset = 1'b0;
	end
	else begin
		case(estado)
			Fetch1: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b1;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Espera1Fetch;
			end
			Espera1Fetch: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b1;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Espera2Fetch;
			end
			Espera2Fetch: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b1;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch2;
			end
			Fetch2: begin
				PCWrite = 1'b1;
				MemCtrl = 1'b0;
				IRWrite = 1'b1;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b1;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Decode1;
			end
			Decode1: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b11;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = EsperaDecode;
			end
			EsperaDecode: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b1;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b11;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Decode2;
			end
			Decode2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b1;
				B_Control = 1'b1;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Instrucao;
			end
			Instrucao: begin
				case(OpCode)
					ARIT: begin //aritmeticos
						case(funct)
							ADD: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b01;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b001;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Add2;
							end
							SUB: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b01;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b010;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Sub2;
							end
							AND: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b01;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b011;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = And2;
							end
							BREAK: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b01;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b010;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Break2;
							end
							RTE: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b010;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Rte2;
							end
							SLL: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b10;
								ShiftAmt = 2'b10;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Sll2;
							end
							SLLV: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Sllv2;
							end
							SRL: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b10;
								ShiftAmt = 2'b10;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Srl2;
							end
							SRA: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b10;
								ShiftAmt = 2'b10;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Sra2;
							end
							SRAV: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Srav2;
							end
							SLT: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b01;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b111;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = Slt2;
							end
							JR: begin
								PCWrite = 1'b1;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b0;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b01;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b000;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0000;
								estado = jr2;
							end
							XCHG: begin
								PCWrite = 1'b0;
								MemCtrl = 1'b0;
								IRWrite = 1'b0;
								A_Control = 1'b0;
								B_Control = 1'b0;
								RegControl = 1'b1;
								ALUOutControl = 1'b0;
								EPCWrite = 1'b0;
								MDControl = 1'b0;
								HI_Control = 1'b0;
								LO_Control = 1'b0;
								IorD = 2'b00;
								ALUSrcA = 2'b00;
								ALUSrcB = 2'b00;
								ExcpCtrl = 2'b00;
								ShiftSrc = 2'b00;
								ShiftAmt = 2'b00;
								SSControl = 2'b00;
								LSControl = 2'b00;
								RegDst = 3'b100;
								PCSource = 3'b000;
								ALUControl = 3'b000;
								ShiftControl = 3'b000;
								DataSrc = 4'b0111;
								estado = xchg2;
							end
						endcase
					end
					ADDI: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = Addi2;
					end
					ADDIU: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = Addiu2;
					end
					J: begin
						PCWrite = 1'b1;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b00;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b100;
						ALUControl = 3'b000;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = j2;
					end
					JAL: begin
						PCWrite = 1'b1;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b1;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b00;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b011;
						PCSource = 3'b100;
						ALUControl = 3'b000;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = jal2;
					end
					LUI: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b00;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b01;
						ShiftAmt = 2'b01;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b000;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = lui2;
					end
					SLTI: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b111;
						ShiftControl = 3'b000;
						DataSrc = 4'b0100;
						estado = slti2;
					end
					BEQ: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b111;
						ShiftControl = 3'b000;
						DataSrc = 4'b0100;
						estado = beq2;
					end
					BNE: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b111;
						ShiftControl = 3'b000;
						DataSrc = 4'b0100;
						estado = bne2;
					end
					BLE: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b111;
						ShiftControl = 3'b000;
						DataSrc = 4'b0100;
						estado = ble2;
					end
					BGT: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b111;
						ShiftControl = 3'b000;
						DataSrc = 4'b0100;
						estado = bgt2;
					end
					SB: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b10;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = sb2;
					end
					LB: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b01;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = lb2;
					end
					LW: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b01;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = lw2;
					end
					LH: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b01;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = lh2;
					end
					SH: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b10;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b01;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = sh2;
					end
					SW: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b1;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b10;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b10;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b10;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b001;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = sw2;
					end
					BLM: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b01;
						ALUSrcA = 2'b01;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b10;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b000;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = blm2;
					end
					default: begin
						PCWrite = 1'b0;
						MemCtrl = 1'b0;
						IRWrite = 1'b0;
						A_Control = 1'b0;
						B_Control = 1'b0;
						RegControl = 1'b0;
						ALUOutControl = 1'b0;
						EPCWrite = 1'b0;
						MDControl = 1'b0;
						HI_Control = 1'b0;
						LO_Control = 1'b0;
						IorD = 2'b00;
						ALUSrcA = 2'b00;
						ALUSrcB = 2'b00;
						ExcpCtrl = 2'b00;
						ShiftSrc = 2'b00;
						ShiftAmt = 2'b00;
						SSControl = 2'b00;
						LSControl = 2'b00;
						RegDst = 3'b000;
						PCSource = 3'b000;
						ALUControl = 3'b000;
						ShiftControl = 3'b000;
						DataSrc = 4'b0000;
						estado = INEXISTENTE;
					end
				endcase
			end
			Add2: begin
				if (overflow) begin
					estado = OVERFLOW;
				end
				else begin
					PCWrite = 1'b0;
					MemCtrl = 1'b0;
					IRWrite = 1'b0;
					A_Control = 1'b0;
					B_Control = 1'b0;
					RegControl = 1'b0;
					ALUOutControl = 1'b1;
					EPCWrite = 1'b0;
					MDControl = 1'b0;
					HI_Control = 1'b0;
					LO_Control = 1'b0;
					IorD = 2'b00;
					ALUSrcA = 2'b01;
					ALUSrcB = 2'b00;
					ExcpCtrl = 2'b00;
					ShiftSrc = 2'b00;
					ShiftAmt = 2'b00;
					SSControl = 2'b00;
					LSControl = 2'b00;
					RegDst = 3'b001;
					PCSource = 3'b000;
					ALUControl = 3'b001;
					ShiftControl = 3'b000;
					DataSrc = 4'b0000;
					estado = AddSubAnd;
				end
			end
			Sub2: begin
				if (overflow) begin
					estado = OVERFLOW;
				end
				else begin
					PCWrite = 1'b0;
					MemCtrl = 1'b0;
					IRWrite = 1'b0;
					A_Control = 1'b0;
					B_Control = 1'b0;
					RegControl = 1'b0;
					ALUOutControl = 1'b1;
					EPCWrite = 1'b0;
					MDControl = 1'b0;
					HI_Control = 1'b0;
					LO_Control = 1'b0;
					IorD = 2'b00;
					ALUSrcA = 2'b01;
					ALUSrcB = 2'b00;
					ExcpCtrl = 2'b00;
					ShiftSrc = 2'b00;
					ShiftAmt = 2'b00;
					SSControl = 2'b00;
					LSControl = 2'b00;
					RegDst = 3'b001;
					PCSource = 3'b000;
					ALUControl = 3'b010;
					ShiftControl = 3'b000;
					DataSrc = 4'b0000;
					estado = AddSubAnd;
				end
			end
			And2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b1;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b011;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = AddSubAnd;
			end
			AddSubAnd: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = AddSubAnd2;
			end
			AddSubAnd2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			Addi2: begin
				if (overflow) begin
					estado = OVERFLOW;
				end
				else begin
					PCWrite = 1'b0;
					MemCtrl = 1'b0;
					IRWrite = 1'b0;
					A_Control = 1'b0;
					B_Control = 1'b0;
					RegControl = 1'b0;
					ALUOutControl = 1'b1;
					EPCWrite = 1'b0;
					MDControl = 1'b0;
					HI_Control = 1'b0;
					LO_Control = 1'b0;
					IorD = 2'b00;
					ALUSrcA = 2'b01;
					ALUSrcB = 2'b10;
					ExcpCtrl = 2'b00;
					ShiftSrc = 2'b00;
					ShiftAmt = 2'b00;
					SSControl = 2'b00;
					LSControl = 2'b00;
					RegDst = 3'b000;
					PCSource = 3'b000;
					ALUControl = 3'b001;
					ShiftControl = 3'b000;
					DataSrc = 4'b0000;
					estado = Addi3;
				end
			end
			Addi3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Addi4;
			end
			Addi4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			Break2: begin
				PCWrite = 1'b1;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b010;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Break3;
			end
			Break3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b010;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			Rte2: begin
				PCWrite = 1'b1;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b010;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			Sll2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0000;
				estado = Sll3;
			end
			Sllv2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0000;
				estado = Sllv3;
			end
			Sll3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b010;
				DataSrc = 4'b0101;
				estado = Sll4;
			end
			Sllv3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b010;
				DataSrc = 4'b0101;
				estado = Sll4;
			end
			Sll4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0101;
				estado = Fetch1;
			end
			Srl2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0101;
				estado = Srl3;
			end
			Srl3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b011;
				DataSrc = 4'b0101;
				estado = Sll4;
			end
			Sra2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0101;
				estado = Sra3;
			end
			Sra3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b10;
				ShiftAmt = 2'b10;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b100;
				DataSrc = 4'b0101;
				estado = Sll4;
			end
			Srav2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0000;
				estado = Srav3;
			end
			Srav3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b100;
				DataSrc = 4'b0101;
				estado = Sll4;
			end
			Addiu2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b1;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Addiu3;
			end
			Addiu3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Addi4;
			end
			Slt2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = Slt3;
			end
			Slt3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b001;
				PCSource = 3'b000;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = Fetch1;
			end
			jr2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			xchg2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b100;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0111;
				estado = xchg3;
			end
			xchg3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0110;
				estado = xchg4;
			end
			xchg4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0110;
				estado = Fetch1;
			end
			j2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b100;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			jal2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b011;
				PCSource = 3'b100;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			lui2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b01;
				ShiftAmt = 2'b01;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b001;
				DataSrc = 4'b0000;
				estado = lui3;
			end
			lui3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b01;
				ShiftAmt = 2'b01;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b010;
				DataSrc = 4'b0101;
				estado = lui4;
			end
			lui4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b01;
				ShiftAmt = 2'b01;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0101;
				estado = Fetch1;
			end
			slti2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = slti3;
			end
			slti3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = Fetch1;
			end
			beq2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = beq3;
			end
			beq3: begin
				if (EQF) begin
					PCWrite = 1'b1;
				end
				else begin
					PCWrite = 1'b0;
				end
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = beq4;
			end
			beq4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = Fetch1;
			end
			bne2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = bne3;
			end
			bne3: begin
				if (!EQF) begin
					PCWrite = 1'b1;
				end
				else begin
					PCWrite = 1'b0;
				end
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = beq4;
			end
			ble2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = ble3;
			end
			ble3: begin
				if (!GTF) begin
					PCWrite = 1'b1;
				end
				else begin
					PCWrite = 1'b0;
				end
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = beq4;
			end
			bgt2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = bgt3;
			end
			bgt3: begin
				if (GTF) begin
					PCWrite = 1'b1;
				end
				else begin
					PCWrite = 1'b0;
				end
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b00;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0100;
				estado = beq4;
			end
			OVERFLOW: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b01;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = overflow2;
			end
			overflow2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b01;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = overflow3;
			end
			overflow3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b01;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b011;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = overflow4;
			end
			overflow4: begin
				PCWrite = 1'b1;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b1;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b01;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b011;
				ALUControl = 3'b010;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = overflow5;
			end
			overflow5: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b01;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			sb2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = sbWait;
			end
			sbWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = sbWait2;
			end
			sbWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b1;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = sb3;
			end
			sb3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			lb2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = lbWait;
			end
			lbWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lbWait2;
			end
			lbWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lbWait3;
			end
			lbWait3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lb3;
			end
			lb3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = Fetch1;
			end
			lh2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b01;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = lhWait;
			end
			lhWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b01;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lhWait2;
			end
			lhWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b01;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lhWait3;
			end
			lhWait3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b01;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lh3;
			end
			lh3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b01;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = Fetch1;
			end
			lw2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = lwWait;
			end
			lwWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lwWait2;
			end
			lwWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b1;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lwWait3;
			end
			lwWait3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = lw3;
			end
			lw3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0001;
				estado = Fetch1;
			end
			sh2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b01;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = shWait;
			end
			shWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b01;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = shWait2;
			end
			shWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b1;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b01;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = sh3;
			end
			sh3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b01;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			sw2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b10;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = swWait;
			end
			swWait: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b10;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = swWait2;
			end
			swWait2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b1;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b10;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = sw3;
			end
			sw3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b10;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b10;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b001;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			blm2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b01;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = blm3;
			end
			blm3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b10;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = blm4;
			end
			blm4: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b10;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = blm5;
			end
			blm5: begin
				if (!EQF && !GTF) begin
					PCWrite = 1'b1;
				end
				else begin
					PCWrite = 1'b0;
				end
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b10;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = blm6;
			end
			blm6: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b01;
				ALUSrcA = 2'b10;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b10;
				RegDst = 3'b000;
				PCSource = 3'b001;
				ALUControl = 3'b111;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
			INEXISTENTE: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = inexistente2;
			end
			inexistente2: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = inexistente3;
			end
			inexistente3: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b00;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b011;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = inexistente4;
			end
			inexistente4: begin
				PCWrite = 1'b1;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b1;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b011;
				ALUControl = 3'b010;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = inexistente5;
			end
			inexistente5: begin
				PCWrite = 1'b0;
				MemCtrl = 1'b0;
				IRWrite = 1'b0;
				A_Control = 1'b0;
				B_Control = 1'b0;
				RegControl = 1'b0;
				ALUOutControl = 1'b0;
				EPCWrite = 1'b0;
				MDControl = 1'b0;
				HI_Control = 1'b0;
				LO_Control = 1'b0;
				IorD = 2'b10;
				ALUSrcA = 2'b00;
				ALUSrcB = 2'b01;
				ExcpCtrl = 2'b00;
				ShiftSrc = 2'b00;
				ShiftAmt = 2'b00;
				SSControl = 2'b00;
				LSControl = 2'b00;
				RegDst = 3'b000;
				PCSource = 3'b000;
				ALUControl = 3'b000;
				ShiftControl = 3'b000;
				DataSrc = 4'b0000;
				estado = Fetch1;
			end
		endcase
	end
end

endmodule: Controle